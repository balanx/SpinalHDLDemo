// Generator : SpinalHDL v1.7.2    git head : 08fc866bebdc40c471ebe327bface63e34406489
// Component : Inout_1
// Git hash  : 23d564a3e9d4d768c2cb1641ec7dc2becc0d2602

`timescale 1ns/1ps

module Inout_1 (
);


  ddrCtrl ddrCtrlInst (
    .signal (signal)  //~
  );
  ddrModel ddrModelInst (
    .signal (signal)  //~
  );

endmodule
